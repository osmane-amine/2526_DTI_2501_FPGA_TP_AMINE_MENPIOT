library ieee;
use ieee.std_logic_1164.all;

entity led_blink is
    port (
        i_clk : in std_logic;
        i_rst_n : in std_logic;
        o_led : out std_logic
    );
end entity led_blink;

architecture rtl of led_blink is
    signal r_led : std_logic := '0';
begin
    process(i_clk, i_rst_n)
	 variable counter : natural range 0 to 5000000 := 0;
    begin
        if (i_rst_n = '0') then
            r_led <= '0';
				counter := 0;
        elsif (rising_edge(i_clk)) then
            if (counter = 5000000) then
					counter := 0;
					r_led <= not r_led;
				else
					counter := counter + 1;
				end if;
        end if;
    end process;
    o_led <= r_led;
end architecture rtl;