library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library pll;
use pll.all;

entity telecran is
    port (
        -- FPGA
        i_clk_50: in std_logic;

        -- HDMI
        io_hdmi_i2c_scl       : inout std_logic;
        io_hdmi_i2c_sda       : inout std_logic;
        o_hdmi_tx_clk        : out std_logic;
        o_hdmi_tx_d          : out std_logic_vector(23 downto 0);
        o_hdmi_tx_de         : out std_logic;
        o_hdmi_tx_hs         : out std_logic;
        i_hdmi_tx_int        : in std_logic;
        o_hdmi_tx_vs         : out std_logic;

        -- KEYs
        i_rst_n : in std_logic;
		  
		-- LEDs
--		o_leds : out std_logic_vector(9 downto 0);
--		o_de10_leds : out std_logic_vector(7 downto 0);

		-- Coder
		i_left_ch_a : in std_logic;
		i_left_ch_b : in std_logic;
		i_left_pb : in std_logic;
		i_right_ch_a : in std_logic;
		i_right_ch_b : in std_logic;
		i_right_pb : in std_logic
    );
end entity telecran;

architecture rtl of telecran is

	constant h_res : natural := 720;
    constant v_res : natural := 480;
	constant mem_size : natural := h_res * v_res;
	constant data_width : natural := 8;

	component I2C_HDMI_Config 
		port (
			iCLK : in std_logic;
			iRST_N : in std_logic;
			I2C_SCLK : out std_logic;
			I2C_SDAT : inout std_logic;
			HDMI_TX_INT  : in std_logic
		);
	 end component;
	 
	component pll 
		port (
			refclk : in std_logic;
			rst : in std_logic;
			outclk_0 : out std_logic;
			locked : out std_logic
		);
	end component;

	component hdmi_controler
		port (
			i_clk : in std_logic;
			i_rst_n : in std_logic;
			o_hdmi_hs : out std_logic;
			o_hdmi_vs : out std_logic;
			o_hdmi_de : out std_logic;
			o_pixel_en : out std_logic;
			o_pixel_address : out natural range 0 to (h_res * v_res - 1);
			o_x_counter : out natural range 0 to (h_res - 1);
			o_y_counter : out natural range 0 to (v_res - 1)
		);
	end component;

	component detector
		generic (
			MAX: natural
		);
		port(
			i_clk_50: in std_logic;
			i_rst_n:in std_logic;
			i_en:in std_logic;
			i_ch_a:in std_logic;
			i_ch_b:in std_logic;
			o_count:out natural range 0 to MAX-1;
		);
	end component detector;

	component dpram
		generic (
			mem_size    : natural := 720 * 480;
			data_width  : natural := 8
		);
		port (
			i_clk_a     : in std_logic;
			i_clk_b     : in std_logic;
			i_data_a    : in std_logic_vector(data_width-1 downto 0);
			i_data_b    : in std_logic_vector(data_width-1 downto 0);
			i_addr_a    : in natural range 0 to mem_size-1;
			i_addr_b    : in natural range 0 to mem_size-1;
			i_we_a      : in std_logic;
			i_we_b      : in std_logic;
			o_q_a       : out std_logic_vector(data_width-1 downto 0);
			o_q_b       : out std_logic_vector(data_width-1 downto 0)
		);
	end component dpram;


	signal s_clk_27 : std_logic;
	signal s_rst_n : std_logic;	-- holds reset as long as pll is not locked
	
	signal s_x_counter : natural range 0 to (h_res - 1);
	signal s_y_counter : natural range 0 to (v_res - 1);
	signal s_pixel_address : natural range 0 to (h_res * v_res - 1);
	signal s_pixel_en : std_logic;

	signal s_x_pos : natural range 0 to (h_res - 1);
	signal s_y_pos : natural range 0 to (v_res - 1);

	signal s_pixel_data : std_logic_vector(data_width-1 downto 0);

begin
--	o_leds <= (others => '0');
--	o_de10_leds <= (others => '0');
	
	-- Frequency for HDMI is 27MHz generated by this PLL
	pll0 : component pll 
		port map (
			refclk => i_clk_50,
			rst => not(i_rst_n),
			outclk_0 => s_clk_27,
			locked => s_rst_n
		);
	
	hdmi_controler0 : component hdmi_controler
		port map (
			i_clk => s_clk_27,
			i_rst_n => s_rst_n,
			o_hdmi_hs => o_hdmi_tx_hs,
			o_hdmi_vs => o_hdmi_tx_vs,
			o_hdmi_de => o_hdmi_tx_de,
			o_pixel_en => open,
			o_pixel_address => open,
			o_x_counter => s_x_counter,
			o_y_counter => s_y_counter
		);

	detector_left : component detector
		generic map (
			MAX:= v_res
		);

		port map (
			i_clk_50 => i_clk_50,
			i_rst_n => i_left_pb,
			i_en => '1',
			i_ch_a => i_left_ch_a,
			i_ch_b => i_left_ch_b,
			o_count => s_y_pos
		);

	detector_right : component detector
		generic map (
			MAX:= h_res
		);

		port map (
			i_clk_50 => i_clk_50,
			i_rst_n => i_right_pb,
			i_en => '1',
			i_ch_a => i_right_ch_a,
			i_ch_b => i_right_ch_b,
			o_count => s_x_pos
		);

	dpram0 : component dpram
		generic map (
			mem_size => h_res * v_res,
			data_width => 8
		);
		port map (
			i_clk_a => s_clk_27,
			i_clk_b => s_clk_27,
			i_data_a => (others => '1'),
			i_data_b => (others => '0'),
			i_addr_a => s_x_pos + s_y_pos * v_res,
			i_addr_b => s_x_counter + s_y_counter * v_res,
			i_we_a => '1',
			i_we_b => '0',
			o_q_a => open,
			o_q_b => s_pixel_data 
		);
	
	-- Connect pixel data
	o_hdmi_tx_clk <= s_clk_27;

	-- CONTRÔLEUR HDMI
--	o_hdmi_tx_d(23 downto 16) <= std_logic_vector(to_unsigned(s_x_counter, 8));
--	o_hdmi_tx_d(15 downto 8) <= std_logic_vector(to_unsigned(s_y_counter, 8));
--	o_hdmi_tx_d(7 downto 0) <= (others => '0');

	-- DÉPLACEMENT D'UN PIXEL
--	o_hdmi_tx_d(23 downto 0) <= (others => '1') when (s_x_counter = s_x_pos and s_y_counter = s_y_pos) else (others => '0');

	-- MÉMORISATION
	o_hdmi_tx_d(23 downto 16) <= s_pixel_data(7 downto 0);
	o_hdmi_tx_d(15 downto 8) <= s_pixel_data(7 downto 0);
	o_hdmi_tx_d(7 downto 0) <= s_pixel_data(7 downto 0);


	-- Configures the ADV7513 for 480p
	I2C_HDMI_Config0 : component I2C_HDMI_Config 
		port map (
			iCLK => i_clk_50,
			iRST_N => i_rst_n,
			I2C_SCLK => io_hdmi_i2c_scl,
			I2C_SDAT => io_hdmi_i2c_sda,
			HDMI_TX_INT => i_hdmi_tx_int
	 );
end architecture rtl;
